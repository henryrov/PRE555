magic
tech sky130A
timestamp 1753353008
<< nwell >>
rect 2855 835 3110 925
rect 2855 725 2910 835
rect 2405 170 2830 310
<< nmos >>
rect 2345 1125 2360 2325
rect 2410 1125 2425 2325
rect 2475 1125 2490 2325
rect 2540 1125 2555 2325
rect 2605 1125 2620 2325
rect 2670 1125 2685 2325
<< ndiff >>
rect 2295 1210 2345 2325
rect 2295 1140 2310 1210
rect 2330 1140 2345 1210
rect 2295 1125 2345 1140
rect 2360 2310 2410 2325
rect 2360 2240 2375 2310
rect 2395 2240 2410 2310
rect 2360 1125 2410 2240
rect 2425 1210 2475 2325
rect 2425 1140 2440 1210
rect 2460 1140 2475 1210
rect 2425 1125 2475 1140
rect 2490 2310 2540 2325
rect 2490 2240 2505 2310
rect 2525 2240 2540 2310
rect 2490 1125 2540 2240
rect 2555 1210 2605 2325
rect 2555 1140 2570 1210
rect 2590 1140 2605 1210
rect 2555 1125 2605 1140
rect 2620 2310 2670 2325
rect 2620 2240 2635 2310
rect 2655 2240 2670 2310
rect 2620 1125 2670 2240
rect 2685 1210 2735 2325
rect 2685 1140 2700 1210
rect 2720 1140 2735 1210
rect 2685 1125 2735 1140
<< ndiffc >>
rect 2310 1140 2330 1210
rect 2375 2240 2395 2310
rect 2440 1140 2460 1210
rect 2505 2240 2525 2310
rect 2570 1140 2590 1210
rect 2635 2240 2655 2310
rect 2700 1140 2720 1210
<< poly >>
rect 2345 2325 2360 2340
rect 2410 2325 2425 2340
rect 2475 2325 2490 2340
rect 2540 2325 2555 2340
rect 2605 2325 2620 2340
rect 2670 2325 2685 2340
rect 2345 1110 2360 1125
rect 2410 1110 2425 1125
rect 2475 1110 2490 1125
rect 2540 1110 2555 1125
rect 2605 1110 2620 1125
rect 2670 1110 2685 1125
rect 2345 1100 2685 1110
rect 2345 1080 2355 1100
rect 2675 1080 2685 1100
rect 2345 1070 2685 1080
<< polycont >>
rect 2355 1080 2675 1100
<< locali >>
rect 2365 2310 2665 2320
rect 2365 2240 2375 2310
rect 2655 2240 2665 2310
rect 2365 2230 2665 2240
rect 430 1450 470 1695
rect 430 1430 440 1450
rect 460 1430 470 1450
rect 2240 1445 2755 1485
rect 2715 1435 2755 1445
rect 430 1420 470 1430
rect 2715 1415 2725 1435
rect 2745 1415 2755 1435
rect 2715 1405 2755 1415
rect 2300 1210 2730 1220
rect 2300 1140 2310 1210
rect 2720 1140 2730 1210
rect 2300 1130 2730 1140
rect 2345 1100 2685 1110
rect 2345 1080 2355 1100
rect 2675 1080 2685 1100
rect 2345 1070 2685 1080
rect 430 445 470 835
rect 2260 685 2410 725
rect 2820 685 2905 725
rect 2260 560 2390 685
rect 2805 645 2855 655
rect 2805 625 2815 645
rect 2845 625 2855 645
rect 2805 615 2855 625
rect 2240 520 2390 560
rect 430 425 440 445
rect 460 425 470 445
rect 430 415 470 425
rect 2265 160 2405 170
rect 2530 160 2625 170
rect 2265 140 2275 160
rect 2265 130 2405 140
rect 2530 130 2625 140
<< viali >>
rect 2375 2240 2395 2310
rect 2395 2240 2505 2310
rect 2505 2240 2525 2310
rect 2525 2240 2635 2310
rect 2635 2240 2655 2310
rect 440 1430 460 1450
rect 1725 1430 1775 1450
rect 1875 1430 1925 1450
rect 2725 1415 2745 1435
rect 2310 1140 2330 1210
rect 2330 1140 2440 1210
rect 2440 1140 2460 1210
rect 2460 1140 2570 1210
rect 2570 1140 2590 1210
rect 2590 1140 2700 1210
rect 2700 1140 2720 1210
rect 2355 1080 2675 1100
rect 2725 695 2745 715
rect 3000 695 3020 715
rect 2815 625 2845 645
rect 1725 505 1775 525
rect 1875 505 1925 525
rect 440 425 460 445
rect 2275 140 2460 160
rect 2500 140 2675 160
rect 2720 140 2740 160
<< metal1 >>
rect 0 2495 100 2565
rect 465 2275 610 2495
rect 490 2120 610 2275
rect 775 2320 875 2565
rect 1550 2515 1650 2565
rect 1550 2510 1935 2515
rect 1550 2470 1870 2510
rect 1930 2470 1935 2510
rect 1550 2465 1935 2470
rect 2325 2420 2425 2565
rect 1715 2415 2425 2420
rect 1715 2375 1720 2415
rect 1780 2375 2425 2415
rect 1715 2370 2425 2375
rect 775 2310 2665 2320
rect 775 2240 2375 2310
rect 2655 2240 2665 2310
rect 775 2230 2665 2240
rect 490 1630 3110 2120
rect 2240 1510 3110 1630
rect 430 1455 1785 1460
rect 430 1450 1720 1455
rect 430 1430 440 1450
rect 460 1430 1720 1450
rect 430 1425 1720 1430
rect 1780 1425 1785 1455
rect 430 1420 1785 1425
rect 1865 1455 1935 1460
rect 1865 1425 1870 1455
rect 1930 1425 1935 1455
rect 1865 1420 1935 1425
rect 2715 1440 2755 1445
rect 2715 1410 2720 1440
rect 2750 1410 2755 1440
rect 2715 1405 2755 1410
rect 2225 1210 2730 1220
rect 2225 1140 2310 1210
rect 2720 1140 2730 1210
rect 2225 1125 2730 1140
rect 2345 1105 2685 1110
rect 2345 1075 2350 1105
rect 2680 1075 2685 1105
rect 2345 1070 2685 1075
rect 315 875 2240 985
rect 2905 975 3110 1510
rect 2300 875 3110 975
rect 315 220 415 875
rect 2300 825 2360 875
rect 2905 835 3110 875
rect 490 770 2360 825
rect 490 715 2265 770
rect 2240 590 2265 715
rect 2355 590 2360 770
rect 2715 720 2755 725
rect 2715 690 2720 720
rect 2750 690 2755 720
rect 2715 685 2755 690
rect 2990 720 3030 725
rect 2990 690 2995 720
rect 3025 690 3030 720
rect 2990 685 3030 690
rect 2805 650 2855 655
rect 2805 620 2810 650
rect 2850 620 2855 650
rect 2805 615 2855 620
rect 2240 585 2360 590
rect 1715 530 1785 535
rect 1715 500 1720 530
rect 1780 500 1785 530
rect 1715 495 1785 500
rect 1865 525 1935 535
rect 1865 505 1875 525
rect 1925 505 1935 525
rect 1865 460 1935 505
rect 2905 485 3110 580
rect 430 445 1935 460
rect 430 425 440 445
rect 460 425 1935 445
rect 430 420 1935 425
rect 430 415 470 420
rect 2240 410 3110 485
rect 2260 280 2415 285
rect 2260 200 2265 280
rect 2355 200 2415 280
rect 2260 195 2415 200
rect 2610 195 2625 285
rect 2265 165 2470 170
rect 2265 135 2270 165
rect 2465 135 2470 165
rect 2265 130 2470 135
rect 2490 165 2690 170
rect 2490 135 2495 165
rect 2685 135 2690 165
rect 2490 130 2690 135
rect 2710 165 2750 170
rect 2710 135 2715 165
rect 2745 135 2750 165
rect 2710 130 2750 135
rect 455 60 2405 110
rect 445 20 2405 60
rect 2610 20 2625 110
rect 445 0 2240 20
rect 0 -70 100 0
rect 775 -25 875 -20
rect 775 -65 780 -25
rect 870 -65 875 -25
rect 775 -70 875 -65
rect 1550 -25 1650 -20
rect 1550 -65 1555 -25
rect 1645 -65 1650 -25
rect 1550 -70 1650 -65
rect 2325 -25 2425 -20
rect 2325 -65 2330 -25
rect 2420 -65 2425 -25
rect 2325 -70 2425 -65
<< via1 >>
rect 1870 2470 1930 2510
rect 1720 2375 1780 2415
rect 1720 1450 1780 1455
rect 1720 1430 1725 1450
rect 1725 1430 1775 1450
rect 1775 1430 1780 1450
rect 1720 1425 1780 1430
rect 1870 1450 1930 1455
rect 1870 1430 1875 1450
rect 1875 1430 1925 1450
rect 1925 1430 1930 1450
rect 1870 1425 1930 1430
rect 2720 1435 2750 1440
rect 2720 1415 2725 1435
rect 2725 1415 2745 1435
rect 2745 1415 2750 1435
rect 2720 1410 2750 1415
rect 2350 1100 2680 1105
rect 2350 1080 2355 1100
rect 2355 1080 2675 1100
rect 2675 1080 2680 1100
rect 2350 1075 2680 1080
rect 2265 590 2355 770
rect 2720 715 2750 720
rect 2720 695 2725 715
rect 2725 695 2745 715
rect 2745 695 2750 715
rect 2720 690 2750 695
rect 2995 715 3025 720
rect 2995 695 3000 715
rect 3000 695 3020 715
rect 3020 695 3025 715
rect 2995 690 3025 695
rect 2810 645 2850 650
rect 2810 625 2815 645
rect 2815 625 2845 645
rect 2845 625 2850 645
rect 2810 620 2850 625
rect 1720 525 1780 530
rect 1720 505 1725 525
rect 1725 505 1775 525
rect 1775 505 1780 525
rect 1720 500 1780 505
rect 2265 200 2355 280
rect 2270 160 2465 165
rect 2270 140 2275 160
rect 2275 140 2460 160
rect 2460 140 2465 160
rect 2270 135 2465 140
rect 2495 160 2685 165
rect 2495 140 2500 160
rect 2500 140 2675 160
rect 2675 140 2685 160
rect 2495 135 2685 140
rect 2715 160 2745 165
rect 2715 140 2720 160
rect 2720 140 2740 160
rect 2740 140 2745 160
rect 2715 135 2745 140
rect 780 -65 870 -25
rect 1555 -65 1645 -25
rect 2330 -65 2420 -25
<< metal2 >>
rect 1865 2510 1935 2515
rect 1865 2470 1870 2510
rect 1930 2470 1935 2510
rect 1715 2415 1785 2420
rect 1715 2375 1720 2415
rect 1780 2375 1785 2415
rect 1715 1455 1785 2375
rect 1715 1425 1720 1455
rect 1780 1425 1785 1455
rect 1715 1420 1785 1425
rect 1865 1455 1935 2470
rect 1865 1425 1870 1455
rect 1930 1425 1935 1455
rect 1865 1420 1935 1425
rect 2715 1440 2755 1445
rect 2715 1410 2720 1440
rect 2750 1410 2755 1440
rect 2345 1105 2690 1110
rect 2345 1075 2350 1105
rect 2680 1075 2690 1105
rect 2345 1070 2690 1075
rect 2260 770 2360 775
rect 2260 590 2265 770
rect 2355 590 2360 770
rect 775 530 1785 535
rect 775 500 1720 530
rect 1780 500 1785 530
rect 775 495 1785 500
rect 775 -25 875 495
rect 2260 280 2360 590
rect 2260 200 2265 280
rect 2355 200 2360 280
rect 2260 195 2360 200
rect 775 -65 780 -25
rect 870 -65 875 -25
rect 775 -70 875 -65
rect 1550 165 2470 170
rect 1550 135 2270 165
rect 2465 135 2470 165
rect 1550 130 2470 135
rect 2490 165 2690 1070
rect 2715 720 2755 1410
rect 2715 690 2720 720
rect 2750 690 2755 720
rect 2715 685 2755 690
rect 2990 720 3030 725
rect 2990 690 2995 720
rect 3025 690 3030 720
rect 2490 135 2495 165
rect 2685 135 2690 165
rect 2490 130 2690 135
rect 2710 650 2855 655
rect 2710 620 2810 650
rect 2850 620 2855 650
rect 2710 615 2855 620
rect 2710 165 2850 615
rect 2710 135 2715 165
rect 2745 135 2850 165
rect 2710 130 2850 135
rect 1550 -25 1650 130
rect 2990 -20 3030 690
rect 1550 -65 1555 -25
rect 1645 -65 1650 -25
rect 1550 -70 1650 -65
rect 2325 -25 3030 -20
rect 2325 -65 2330 -25
rect 2420 -65 3030 -25
rect 2325 -70 3030 -65
use comp  comp_0
timestamp 1753284924
transform 1 0 550 0 1 0
box -60 0 1690 775
use comp  comp_1
timestamp 1753284924
transform 1 0 550 0 1 925
box -60 0 1690 775
use inverter  inverter_0
timestamp 1753284924
transform -1 0 2710 0 1 35
box -120 -35 85 275
use inverter  inverter_1
timestamp 1753284924
transform -1 0 2490 0 1 35
box -120 -35 85 275
use inverter  inverter_2
timestamp 1753284924
transform -1 0 2990 0 1 590
box -120 -35 85 275
use sr_latch  sr_latch_0
timestamp 1753106794
transform 1 0 2450 0 1 570
box -45 -115 405 355
use vdiv  vdiv_0
timestamp 1753016921
transform 1 0 0 0 1 0
box 0 0 470 2495
<< labels >>
rlabel metal1 0 -70 100 -70 5 GND
port 1 s
rlabel metal1 775 -70 875 -70 5 TRIGGER
port 2 s
rlabel metal1 1550 -70 1650 -70 5 OUTPUT
port 3 s
rlabel metal1 2325 -70 2425 -70 5 RESET
port 4 s
rlabel metal1 0 2565 100 2565 1 VDD
port 5 n
rlabel metal1 775 2565 875 2565 1 DISCHARGE
port 6 n
rlabel metal1 1550 2565 1650 2565 1 THRESHOLD
port 7 n
rlabel metal1 2325 2565 2425 2565 1 CONTROL
port 8 n
<< end >>
