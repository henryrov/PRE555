** sch_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/comp.sch
**.subckt comp inp inn out
*.ipin inp
*.ipin inn
*.opin out
XM1 net1 inn net3 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM2 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM3 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM4 net2 inp net3 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM5 net3 net4 GND GND sky130_fd_pr__nfet_01v8 L=1 W=3.5 nf=1 ad=1.015 as=1.015 pd=7.58 ps=7.58 nrd=0.0828571428571429
+ nrs=0.0828571428571429 sa=0 sb=0 sd=0 mult=1 m=1
XM6 net4 net4 GND GND sky130_fd_pr__nfet_01v8 L=1 W=3.5 nf=1 ad=1.015 as=1.015 pd=7.58 ps=7.58 nrd=0.0828571428571429
+ nrs=0.0828571428571429 sa=0 sb=0 sd=0 mult=1 m=1
XR1 net4 VDD res100k
X1 net2 out inverter
**.ends

* expanding   symbol:  res100k.sym # of pins=2
** sym_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/res100k.sym
** sch_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/res100k.sch
.subckt res100k bot top
*.iopin top
*.iopin bot
XR1 net1 top GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
XR2 net2 net1 GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
XR3 net3 net2 GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
XR4 net4 net3 GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
XR5 bot net4 GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=2
** sym_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/inverter.sym
** sch_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/inverter.sch
.subckt inverter a y
*.ipin a
*.opin y
XM1 y a GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM2 y a VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
