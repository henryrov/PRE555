* NGSPICE file created from comp.ext - technology: sky130A

.subckt inverter a y VDD GND
X0 y a VDD VDD sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 y a GND GND sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

.subckt res100k bot top GND
X0 a_0_668# bot GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X1 top a_348_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X2 a_0_668# a_116_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X3 a_232_668# a_116_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X4 a_232_668# a_348_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
.ends

*.subckt comp inn inp
Xinverter_0 inverter_0/a inverter_0/y VDD GND inverter
Xres100k_0 res100k_0/bot VDD GND res100k
X0 VDD a_2200_760# a_2200_760# VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X1 GND res100k_0/bot a_1460_170# GND sky130_fd_pr__nfet_01v8 ad=3.5 pd=9 as=3.5 ps=9 w=3.5 l=1
X2 inverter_0/a a_2200_760# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
X3 GND res100k_0/bot res100k_0/bot GND sky130_fd_pr__nfet_01v8 ad=3.5 pd=9 as=3.5 ps=9 w=3.5 l=1
X4 a_1460_170# inn a_2200_760# GND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X5 inverter_0/a inp a_1460_170# GND sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
*.ends

