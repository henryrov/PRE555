** sch_path: /home/henryrovner/Repos/ic_design/PRE555/xschem/inverter.sch
**.subckt inverter a y
*.ipin a
*.opin y
XM1 y a GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM2 y a VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
