* SPICE3 file created from inverter.ext - technology: sky130A

*.subckt inverter a y
X0 y a VDD VDD sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 y a GND GND sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
*.ends

