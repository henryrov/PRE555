magic
tech sky130A
timestamp 1753284924
<< nwell >>
rect 1080 675 1690 775
rect 1080 560 1485 675
<< nmos >>
rect 500 85 600 435
rect 830 85 930 435
rect 1150 380 1250 480
rect 1300 380 1400 480
<< pmos >>
rect 1150 595 1250 695
rect 1300 595 1400 695
<< ndiff >>
rect 1100 465 1150 480
rect 400 420 500 435
rect 400 100 415 420
rect 485 100 500 420
rect 400 85 500 100
rect 600 420 700 435
rect 600 100 615 420
rect 685 100 700 420
rect 600 85 700 100
rect 730 420 830 435
rect 730 100 745 420
rect 815 100 830 420
rect 730 85 830 100
rect 930 420 1030 435
rect 930 100 945 420
rect 1015 100 1030 420
rect 1100 395 1115 465
rect 1135 395 1150 465
rect 1100 380 1150 395
rect 1250 465 1300 480
rect 1250 395 1265 465
rect 1285 395 1300 465
rect 1250 380 1300 395
rect 1400 465 1450 480
rect 1400 395 1415 465
rect 1435 395 1450 465
rect 1400 380 1450 395
rect 930 85 1030 100
<< pdiff >>
rect 1100 680 1150 695
rect 1100 610 1115 680
rect 1135 610 1150 680
rect 1100 595 1150 610
rect 1250 680 1300 695
rect 1250 610 1265 680
rect 1285 610 1300 680
rect 1250 595 1300 610
rect 1400 680 1450 695
rect 1400 610 1415 680
rect 1435 610 1450 680
rect 1400 595 1450 610
<< ndiffc >>
rect 415 100 485 420
rect 615 100 685 420
rect 745 100 815 420
rect 945 100 1015 420
rect 1115 395 1135 465
rect 1265 395 1285 465
rect 1415 395 1435 465
<< pdiffc >>
rect 1115 610 1135 680
rect 1265 610 1285 680
rect 1415 610 1435 680
<< psubdiff >>
rect 1075 280 1660 295
rect 1075 20 1090 280
rect 1645 20 1660 280
rect 1075 5 1660 20
<< nsubdiff >>
rect 1245 750 1450 755
rect 1245 730 1260 750
rect 1435 730 1450 750
rect 1245 725 1450 730
<< psubdiffcont >>
rect 1090 20 1645 280
<< nsubdiffcont >>
rect 1260 730 1435 750
<< poly >>
rect 1150 740 1190 750
rect 1150 720 1160 740
rect 1180 720 1190 740
rect 1150 710 1190 720
rect 1150 695 1250 710
rect 1300 695 1400 710
rect 1150 580 1250 595
rect 1300 580 1400 595
rect 1150 560 1400 580
rect 1165 525 1235 535
rect 500 510 930 520
rect 500 460 510 510
rect 590 460 930 510
rect 1165 505 1175 525
rect 1225 505 1235 525
rect 1165 495 1235 505
rect 1315 525 1385 535
rect 1315 505 1325 525
rect 1375 505 1385 525
rect 1315 495 1385 505
rect 1150 480 1250 495
rect 1300 480 1400 495
rect 500 450 930 460
rect 500 435 600 450
rect 830 435 930 450
rect 1150 365 1250 380
rect 1300 365 1400 380
rect 500 70 600 85
rect 830 70 930 85
<< polycont >>
rect 1160 720 1180 740
rect 510 460 590 510
rect 1175 505 1225 525
rect 1325 505 1375 525
<< locali >>
rect -60 765 -20 775
rect -60 725 -50 765
rect -30 725 -20 765
rect -60 220 -20 725
rect 232 555 495 775
rect 1245 750 1450 755
rect 232 554 375 555
rect 405 520 495 555
rect 1105 740 1190 750
rect 1105 720 1160 740
rect 1180 720 1190 740
rect 1245 730 1260 750
rect 1435 730 1450 750
rect 1245 725 1450 730
rect 1105 710 1190 720
rect 1105 680 1145 710
rect 1105 610 1115 680
rect 1135 610 1145 680
rect 405 510 600 520
rect 405 460 510 510
rect 590 460 600 510
rect 405 450 600 460
rect 735 450 1085 520
rect 405 420 495 450
rect -60 0 35 220
rect 330 65 365 350
rect 405 100 415 420
rect 485 100 495 420
rect 405 90 495 100
rect 605 420 695 430
rect 605 100 615 420
rect 685 100 695 420
rect 605 65 695 100
rect 735 420 825 450
rect 735 100 745 420
rect 815 100 825 420
rect 735 90 825 100
rect 935 420 1025 430
rect 935 100 945 420
rect 1015 100 1025 420
rect 1045 360 1085 450
rect 1105 465 1145 610
rect 1255 680 1295 725
rect 1255 610 1265 680
rect 1285 610 1295 680
rect 1255 600 1295 610
rect 1405 680 1445 690
rect 1405 610 1415 680
rect 1435 610 1445 680
rect 1405 560 1445 610
rect 1165 525 1235 535
rect 1165 505 1175 525
rect 1225 505 1235 525
rect 1165 495 1235 505
rect 1315 525 1385 535
rect 1315 505 1325 525
rect 1375 505 1385 525
rect 1315 495 1385 505
rect 1405 520 1570 560
rect 1105 395 1115 465
rect 1135 395 1145 465
rect 1105 385 1145 395
rect 1255 465 1295 475
rect 1255 395 1265 465
rect 1285 395 1295 465
rect 1255 360 1295 395
rect 1405 465 1445 520
rect 1405 395 1415 465
rect 1435 395 1445 465
rect 1405 385 1445 395
rect 1045 320 1295 360
rect 935 65 1025 100
rect 1075 280 1660 295
rect 1075 65 1090 280
rect 330 20 1090 65
rect 1645 20 1660 280
rect 330 5 1660 20
<< viali >>
rect -50 725 -30 765
rect 1260 730 1435 750
rect 1090 20 1645 280
<< metal1 >>
rect -60 765 1690 775
rect -60 725 -50 765
rect -30 750 1690 765
rect -30 730 1260 750
rect 1435 730 1690 750
rect -30 725 1690 730
rect -60 715 1690 725
rect 1485 675 1690 715
rect 1485 295 1690 430
rect 1075 280 1690 295
rect 1075 60 1090 280
rect -60 20 1090 60
rect 1645 20 1690 280
rect -60 0 1690 20
use inverter  inverter_0
timestamp 1753284924
transform 1 0 1605 0 1 425
box -120 -35 85 275
use res100k  res100k_0
timestamp 1753015857
transform -1 0 267 0 -1 554
box -105 -220 267 554
<< labels >>
rlabel metal1 -60 715 1690 775 1 VDD
rlabel metal1 -60 0 1690 60 5 GND
rlabel locali 1165 495 1235 535 1 inn
port 1 n
rlabel locali 1315 495 1385 535 1 inp
port 2 n
rlabel space 1690 520 1690 560 3 out
<< end >>
