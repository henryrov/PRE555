magic
tech sky130A
timestamp 1753106794
<< nwell >>
rect -45 155 405 355
<< nmos >>
rect 0 -55 15 45
rect 55 -55 70 45
rect 225 -55 240 45
rect 280 -55 295 45
rect 335 -55 350 45
<< pmos >>
rect 15 175 30 275
rect 55 175 70 275
rect 225 175 240 275
rect 265 175 280 275
rect 330 175 345 275
<< ndiff >>
rect -40 30 0 45
rect -40 -40 -30 30
rect -10 -40 0 30
rect -40 -55 0 -40
rect 15 30 55 45
rect 15 -40 25 30
rect 45 -40 55 30
rect 15 -55 55 -40
rect 70 30 110 45
rect 70 -40 80 30
rect 100 -40 110 30
rect 70 -55 110 -40
rect 185 30 225 45
rect 185 -40 195 30
rect 215 -40 225 30
rect 185 -55 225 -40
rect 240 30 280 45
rect 240 -40 250 30
rect 270 -40 280 30
rect 240 -55 280 -40
rect 295 30 335 45
rect 295 -40 305 30
rect 325 -40 335 30
rect 295 -55 335 -40
rect 350 30 390 45
rect 350 -40 360 30
rect 380 -40 390 30
rect 350 -55 390 -40
<< pdiff >>
rect -25 260 15 275
rect -25 190 -15 260
rect 5 190 15 260
rect -25 175 15 190
rect 30 175 55 275
rect 70 260 110 275
rect 70 190 80 260
rect 100 190 110 260
rect 70 175 110 190
rect 185 260 225 275
rect 185 190 195 260
rect 215 190 225 260
rect 185 175 225 190
rect 240 175 265 275
rect 280 175 330 275
rect 345 260 385 275
rect 345 190 355 260
rect 375 190 385 260
rect 345 175 385 190
<< ndiffc >>
rect -30 -40 -10 30
rect 25 -40 45 30
rect 80 -40 100 30
rect 195 -40 215 30
rect 250 -40 270 30
rect 305 -40 325 30
rect 360 -40 380 30
<< pdiffc >>
rect -15 190 5 260
rect 80 190 100 260
rect 195 190 215 260
rect 355 190 375 260
<< psubdiff >>
rect -40 -90 390 -85
rect -40 -110 -25 -90
rect 375 -110 390 -90
rect -40 -115 390 -110
<< nsubdiff >>
rect -25 330 385 335
rect -25 310 -10 330
rect 370 310 385 330
rect -25 305 385 310
<< psubdiffcont >>
rect -25 -110 375 -90
<< nsubdiffcont >>
rect -10 310 370 330
<< poly >>
rect 15 275 30 290
rect 55 275 70 290
rect 225 275 240 290
rect 265 275 280 290
rect 330 275 345 290
rect 15 155 30 175
rect -40 145 30 155
rect -40 125 -30 145
rect -10 130 30 145
rect -10 125 15 130
rect -40 115 15 125
rect 0 45 15 115
rect 55 90 70 175
rect 95 145 135 155
rect 225 145 240 175
rect 95 125 105 145
rect 125 125 240 145
rect 95 115 135 125
rect 160 90 200 100
rect 55 70 170 90
rect 190 70 200 90
rect 55 45 70 70
rect 160 60 200 70
rect 225 45 240 125
rect 265 155 280 175
rect 330 155 345 175
rect 265 145 305 155
rect 265 125 275 145
rect 295 125 305 145
rect 265 115 305 125
rect 330 145 370 155
rect 330 125 340 145
rect 360 125 370 145
rect 330 115 370 125
rect 265 70 280 115
rect 330 75 345 115
rect 265 55 295 70
rect 330 60 350 75
rect 280 45 295 55
rect 335 45 350 60
rect 0 -70 15 -55
rect 55 -70 70 -55
rect 225 -70 240 -55
rect 280 -70 295 -55
rect 335 -70 350 -55
<< polycont >>
rect -30 125 -10 145
rect 105 125 125 145
rect 170 70 190 90
rect 275 125 295 145
rect 340 125 360 145
<< locali >>
rect -25 330 385 335
rect -25 310 -10 330
rect 370 310 385 330
rect -25 305 385 310
rect -20 260 10 305
rect -20 190 -15 260
rect 5 190 10 260
rect -20 180 10 190
rect 75 260 105 270
rect 75 190 80 260
rect 100 190 105 260
rect 75 155 105 190
rect 190 260 220 275
rect 190 190 195 260
rect 215 190 220 260
rect -40 145 0 155
rect -40 125 -30 145
rect -10 125 0 145
rect -40 115 0 125
rect 20 145 135 155
rect 20 125 105 145
rect 125 125 135 145
rect 20 115 135 125
rect -35 30 -5 40
rect -35 -40 -30 30
rect -10 -40 -5 30
rect -35 -85 -5 -40
rect 20 30 50 115
rect 190 100 220 190
rect 350 260 380 305
rect 350 190 355 260
rect 375 190 380 260
rect 350 175 380 190
rect 265 145 305 155
rect 265 125 275 145
rect 295 125 305 145
rect 265 115 305 125
rect 330 145 370 155
rect 330 125 340 145
rect 360 125 370 145
rect 330 115 370 125
rect 160 90 220 100
rect 160 70 170 90
rect 190 80 220 90
rect 190 70 405 80
rect 160 60 405 70
rect 20 -40 25 30
rect 45 -40 50 30
rect 20 -50 50 -40
rect 75 30 105 40
rect 75 -40 80 30
rect 100 -40 105 30
rect 75 -85 105 -40
rect 190 30 220 40
rect 190 -40 195 30
rect 215 -40 220 30
rect 190 -85 220 -40
rect 245 30 275 60
rect 245 -40 250 30
rect 270 -40 275 30
rect 245 -50 275 -40
rect 300 30 330 40
rect 300 -40 305 30
rect 325 -40 330 30
rect 300 -85 330 -40
rect 355 30 385 60
rect 355 -40 360 30
rect 380 -40 385 30
rect 355 -50 385 -40
rect -40 -90 390 -85
rect -40 -110 -25 -90
rect 375 -110 390 -90
rect -40 -115 390 -110
<< viali >>
rect -10 310 370 330
rect -25 -110 375 -90
<< metal1 >>
rect -45 330 405 335
rect -45 310 -10 330
rect 370 310 405 330
rect -45 305 405 310
rect -45 -90 405 -85
rect -45 -110 -25 -90
rect 375 -110 405 -90
rect -45 -115 405 -110
<< labels >>
rlabel locali -40 115 0 155 7 s
port 1 w
rlabel locali 405 60 405 80 3 q
port 4 e
rlabel locali 265 115 305 155 7 r0
port 2 w
rlabel locali 330 115 370 155 3 r1
port 3 e
rlabel metal1 -45 305 370 335 1 VDD
rlabel metal1 -45 -115 370 -85 5 GND
<< end >>
