* SPICE3 file created from vdiv.ext - technology: sky130A

.subckt res100k bot top GND
X0 a_0_668# bot GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X1 top a_348_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X2 a_0_668# a_116_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X3 a_232_668# a_116_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X4 a_232_668# a_348_n440# GND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
.ends

*.subckt vdiv v1t v2t
Xres100k_0[0] GND v1t GND res100k
Xres100k_0[1] v1t v2t GND res100k
Xres100k_0[2] v2t VDD GND res100k
*.ends

